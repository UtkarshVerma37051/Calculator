`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:05:17 02/14/2020 
// Design Name: 
// Module Name:    Final_Mul 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Final_Mul(output [7:0] out,input [7:0] A,B,input Sign_A,Sign_B,Rst);
wire [7:0] wa;
wire [7:0] wb;
wire [15:0] s;
Sign_Sel sa(wa[7:0],A[7:0],Sign_A,Rst);
Sign_Sel sb(wb[7:0],B[7:0],Sign_B,Rst);
Mul_8_Bit M0(s[15:0],wa[7:0],wb[7:0],Rst);
assign out[7:0] = s[7:0];

endmodule
